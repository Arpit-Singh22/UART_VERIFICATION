`include "../rtl/uvm_top.v"
`include "../wb_intf/wb_intf.sv"
`include "../top/top.sv"
