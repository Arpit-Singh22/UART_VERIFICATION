typedef uvm_sequencer#(wb_tx) uart_sqr;
