`include "../wb_intf/wb_intf.sv"
`include "../rtl/uart_top.v"
`include "../top/top.sv"
