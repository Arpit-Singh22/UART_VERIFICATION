`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "./uart_controller/uart_controller.sv"

`include "apb_common.sv"
`include "apb_if.sv"

`include "apb_tx.sv"
`include "apb_sequence.sv"
`include "apb_sqr.sv"
`include "apb_driver.sv"
//`include "apb_mon.sv"
//`include "apb_cov.sv"
`include "apb_agent.sv"
`include "apb_env.sv"
`include "apb_test.sv"
`include "top.sv"
